library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.constants.all;

entity main is
	generic(
        COST_W : integer := CONST_COST_W - 1;
        DATA_W : integer := CONST_DATA_W - 1;
        COOR_W : integer := CONST_COOR_W - 1;
        ADDR_W : integer := CONST_ADDR_W - 1
    );
end main;

architecture arquitectura of main is
   component processor_buffer is
        port(
            clk          : in std_logic;
            rst          : in std_logic;
            adv          : in std_logic;
            wrena_l      : in std_logic;
            wrena_r      : in std_logic;
            left         : in std_logic_vector(DATA_W downto 0);
            right        : in std_logic_vector(DATA_W downto 0);
            row          : in std_logic_vector(COOR_W downto 0);
            cost         : out std_logic_vector(COST_W downto 0);
            process_wait : out std_logic
        );
    end component;
    
    component addr_generator is
        port(
            clk        : in std_logic;
            rst        : in std_logic;
            adv        : in std_logic;
            vs         : out std_logic;
            column     : out std_logic_vector(COOR_W downto 0);
            row        : out std_logic_vector(COOR_W downto 0);
            addr_left  : out std_logic_vector(ADDR_W downto 0);
            addr_right : out std_logic_vector(ADDR_W downto 0);
            addr_out   : out std_logic_vector(ADDR_W downto 0)
        );
    end component;
	
	type ARRAY_IMAGE is array (0 to 80) of integer range 0 to 255;
	
	signal i : std_logic_vector(7 downto 0) := (others => '0');
	signal element : std_logic_vector(15 downto 0) := (others => '0');
	
	signal clk : std_logic := '0';
	signal rst : std_logic := '0';
	signal adv : std_logic := '1';
	
    signal counter : std_logic_vector(COOR_W downto 0) := (others => '0');
	signal state   : std_logic_vector(1 downto 0) := b"11";
	signal activate : std_logic_vector(2 downto 0) := (others => '0');
    
    signal in_acumulator  : std_logic_vector(COST_W downto 0); 
	signal out_acumulator : std_logic_vector(COST_W downto 0);	
	signal acumulated     : std_logic_vector(COST_W downto 0);
	
	signal addr_left : std_logic_vector(15 downto 0);
	signal addr_right : std_logic_vector(15 downto 0);
	signal addr_out : std_logic_vector(15 downto 0); 

	signal pixel_left  : std_logic_vector(DATA_W downto 0);
    signal pixel_right : std_logic_vector(DATA_W downto 0);
	

	type t_array_image is array (0 to 3839) of integer range 0 to 255;
	
	
	-- Arreglo que contiene informacion.
	constant buffer_left : t_array_image:= (
		17, 7, 6, 6, 6, 7, 6, 7, 6, 6, 7, 8, 10, 9, 12, 10, 12, 12, 14, 19, 24, 24, 20, 20, 32, 42, 46, 46, 46, 45, 47, 44, 46, 47, 52, 55, 65, 56, 54, 63, 44, 10, 17, 19, 18, 8, 8, 10, 9, 7, 9, 8, 7, 10, 36, 58, 55, 56, 57, 55, 56, 57, 56, 56, 56, 54, 54, 54, 53, 54, 56, 54, 55, 54, 56, 55, 55, 54, 54, 54, 55, 54, 55, 56, 54, 55, 55, 54, 55, 55, 54, 54, 55, 57, 79, 88, 84, 84, 86, 85, 85, 85, 86, 84, 84, 85, 85, 85, 87, 90, 94, 93, 95, 90, 75, 77, 83, 96, 76, 72, 84, 101, 91, 81, 92, 86, 83, 87, 89, 89, 81, 92, 89, 90, 97, 103, 96, 97, 98, 96, 62, 76, 92, 89, 57, 74, 97, 77, 67, 72, 90, 84, 89, 87, 60, 26, 43, 73, 94, 83, 86, 88, 85, 66, 47, 56, 53, 51, 54, 53, 53, 52, 52, 50, 52, 51, 52, 50, 51, 50, 49, 48, 49, 48, 47, 48, 49, 48, 48, 47, 45, 20, 19, 17, 6, 2, 5, 5, 5, 6, 11, 17, 18, 19, 20, 21, 29, 45, 53, 51, 53, 50, 51, 50, 51, 47, 20, 4, 16, 4, 6, 4, 4, 8, 22, 37, 31, 21, 19, 17, 17, 16, 17, 15, 15, 15, 16, 16, 16, 16, 15, 13, 16, 15, 15, 15, 15, 15, 17, 25, 37, 43, 45, 44, 42, 43, 43, 42, 42, 38, 39, 36, 31, 25, 22, 18, 16, 14, 15, 13, 14, 12, 12, 9, 6, 5, 4, 4, 4, 3, 4, 4, 7, 18, 28, 31, 35, 34, 35, 35, 35, 34, 33, 32, 34, 34, 35, 34, 35, 34, 34, 35, 36, 32, 32, 27, 20, 30, 26, 23, 25, 35, 35, 36, 35, 35, 36, 35, 38, 38,
		39, 36, 38, 37, 38, 38, 39, 37, 38, 38, 38, 37, 39, 37, 33, 22, 21, 20, 21, 21, 22, 21, 22, 22, 23, 22, 23, 21, 23, 22, 23, 22, 22, 22, 23, 23, 23, 27, 37, 43, 48, 47, 49, 48, 49, 48, 49, 50, 49, 49, 49, 48, 47, 44, 43, 41, 43, 41, 41, 40, 42, 44, 43, 22, 31, 15, 10, 13, 13, 13, 14, 13, 13, 15, 14, 14, 18, 19, 22, 22, 24, 23, 24, 27, 33, 35, 35, 36, 52, 66, 73, 71, 71, 70, 72, 69, 69, 70, 79, 87, 126, 125, 75, 118, 94, 6, 41, 46, 43, 20, 23, 32, 24, 14, 20, 18, 17, 15, 70, 115, 111, 112, 116, 110, 111, 112, 114, 112, 112, 109, 109, 107, 108, 107, 112, 110, 112, 112, 112, 110, 111, 109, 107, 108, 111, 109, 112, 112, 110, 109, 111, 110, 109, 108, 110, 108, 111, 113, 157, 180, 170, 170, 174, 171, 172, 172, 173, 171, 171, 173, 172, 173, 175, 182, 190, 190, 191, 187, 123, 87, 118, 191, 170, 160, 173, 201, 179, 160, 180, 189, 168, 173, 194, 174, 158, 164, 189, 178, 197, 201, 201, 190, 193, 195, 137, 80, 171, 190, 107, 123, 201, 150, 89, 119, 185, 171, 178, 172, 141, 93, 147, 155, 184, 170, 173, 175, 172, 133, 95, 112, 104, 104, 106, 108, 106, 106, 108, 104, 106, 105, 104, 104, 104, 101, 99, 98, 99, 99, 98, 96, 96, 94, 97, 95, 94, 43, 36, 37, 15, 6, 12, 10, 10, 11, 24, 37, 39, 39, 40, 40, 57, 90, 103, 101, 103, 101, 101, 100, 101, 92, 40, 5, 20, 13, 12, 10, 10, 17, 45, 78, 64, 43, 36, 33, 33, 33, 33, 30, 32, 31, 35, 32, 33, 32, 32, 31, 34, 31, 32, 31, 33, 30, 36, 50, 74, 85, 91, 90, 88, 85,
		85, 84, 83, 77, 75, 66, 55, 45, 40, 33, 32, 29, 29, 28, 29, 26, 26, 20, 13, 11, 11, 8, 9, 8, 9, 9, 16, 37, 56, 63, 71, 68, 71, 69, 70, 69, 66, 62, 70, 68, 70, 69, 69, 68, 68, 69, 72, 66, 66, 54, 42, 60, 54, 47, 51, 71, 71, 73, 71, 71, 73, 72, 77, 77, 77, 76, 77, 75, 77, 78, 78, 76, 78, 78, 77, 77, 77, 76, 65, 44, 44, 44, 44, 43, 45, 44, 43, 45, 46, 45, 47, 47, 45, 45, 46, 45, 46, 46, 46, 46, 48, 56, 75, 88, 94, 93, 93, 94, 97, 95, 98, 96, 94, 96, 96, 93, 93, 89, 87, 86, 88, 86, 85, 81, 81, 81, 79, 39, 27, 15, 11, 15, 13, 13, 13, 13, 13, 13, 14, 14, 18, 20, 22, 20, 23, 23, 23, 24, 28, 29, 31, 33, 42, 50, 52, 48, 46, 44, 43, 39, 37, 33, 35, 37, 43, 48, 46, 50, 52, 35, 49, 52, 46, 20, 19, 52, 46, 9, 19, 19, 17, 16, 63, 112, 109, 111, 112, 109, 113, 112, 111, 111, 110, 108, 109, 108, 112, 110, 112, 109, 112, 111, 114, 110, 111, 110, 109, 107, 110, 110, 110, 110, 112, 112, 112, 107, 109, 109, 109, 106, 111, 113, 153, 178, 168, 169, 173, 171, 173, 171, 174, 171, 171, 170, 173, 173, 176, 182, 190, 190, 191, 188, 155, 99, 120, 176, 186, 152, 176, 204, 180, 156, 175, 194, 176, 179, 193, 171, 159, 176, 189, 176, 195, 199, 210, 194, 190, 195, 135, 103, 175, 180, 103, 129, 200, 147, 99, 127, 187, 167, 179, 172, 118, 107, 111, 144, 191, 165, 177, 174, 171, 135, 94, 110, 105, 104, 107, 105, 106, 105, 107, 107, 106, 105, 105, 104, 105, 101, 99, 97, 99, 98, 98, 96, 97, 95, 98, 97, 93, 45,
		36, 37, 17, 5, 11, 10, 10, 12, 24, 35, 37, 36, 38, 40, 63, 94, 102, 99, 101, 98, 99, 98, 101, 90, 42, 5, 20, 15, 13, 10, 11, 17, 44, 76, 67, 45, 37, 33, 35, 35, 33, 31, 32, 34, 33, 32, 32, 31, 31, 31, 33, 31, 32, 34, 33, 32, 34, 49, 74, 85, 90, 89, 88, 83, 84, 86, 84, 72, 64, 54, 46, 39, 34, 30, 31, 28, 30, 29, 29, 27, 27, 19, 12, 10, 9, 7, 9, 8, 10, 10, 15, 36, 55, 63, 73, 70, 72, 68, 71, 69, 69, 66, 70, 68, 69, 68, 70, 69, 69, 70, 71, 68, 65, 56, 43, 60, 53, 45, 51, 69, 73, 73, 71, 71, 73, 71, 78, 77, 77, 75, 77, 75, 77, 77, 79, 76, 76, 78, 76, 76, 75, 74, 65, 44, 45, 44, 46, 45, 47, 45, 45, 45, 47, 44, 47, 47, 47, 45, 45, 45, 47, 46, 48, 46, 48, 55, 71, 80, 85, 83, 88, 85, 86, 86, 88, 85, 87, 84, 84, 82, 84, 81, 80, 80, 80, 78, 75, 71, 70, 66, 66, 32, 25, 16, 11, 14, 14, 13, 14, 13, 12, 14, 13, 14, 20, 19, 21, 20, 23, 22, 24, 24, 25, 25, 26, 27, 33, 36, 37, 35, 32, 30, 29, 27, 28, 27, 26, 28, 31, 33, 39, 42, 48, 51, 55, 55, 46, 17, 21, 28, 38, 14, 20, 17, 19, 16, 58, 112, 110, 111, 110, 110, 112, 110, 110, 109, 111, 110, 110, 107, 109, 108, 111, 108, 108, 107, 111, 108, 108, 109, 112, 111, 111, 110, 109, 108, 110, 109, 109, 108, 110, 109, 110, 108, 111, 109, 147, 182, 168, 168, 173, 169, 174, 171, 171, 169, 172, 170, 173, 172, 175, 182, 193, 189, 188, 183, 145, 113, 144, 195, 173, 157, 178, 202, 187, 168, 177, 195, 166, 154,
		188, 160, 176, 164, 191, 177, 194, 196, 207, 198, 189, 193, 179, 139, 154, 201, 135, 109, 202, 144, 120, 148, 184, 168, 178, 173, 135, 114, 103, 157, 183, 172, 172, 174, 172, 133, 94, 112, 108, 105, 107, 105, 106, 104, 106, 106, 105, 104, 106, 103, 107, 103, 100, 98, 99, 100, 100, 97, 98, 96, 99, 96, 91, 45, 36, 38, 19, 5, 11, 12, 9, 10, 17, 22, 23, 23, 24, 25, 38, 54, 59, 59, 57, 57, 58, 55, 57, 50, 25, 10, 15, 12, 12, 10, 11, 18, 43, 73, 65, 41, 36, 34, 35, 34, 33, 33, 33, 31, 33, 33, 33, 32, 33, 33, 33, 33, 34, 33, 36, 32, 35, 49, 73, 85, 89, 87, 88, 86, 85, 84, 79, 64, 54, 44, 39, 32, 32, 29, 30, 27, 30, 28, 31, 26, 25, 20, 12, 10, 10, 7, 10, 7, 9, 9, 15, 33, 53, 63, 73, 69, 72, 68, 70, 68, 70, 67, 68, 69, 71, 69, 70, 68, 69, 69, 73, 67, 68, 57, 42, 61, 53, 45, 49, 69, 72, 72, 71, 70, 73, 73, 77, 77, 75, 76, 78, 75, 76, 77, 78, 76, 77, 75, 77, 74, 76, 74, 66, 45, 48, 46, 47, 46, 47, 46, 48, 45, 48, 45, 47, 46, 48, 46, 47, 45, 46, 45, 47, 47, 49, 51, 64, 67, 71, 71, 72, 71, 72, 70, 71, 71, 71, 69, 71, 70, 70, 67, 67, 67, 67, 62, 63, 61, 59, 58, 56, 27, 23, 16, 10, 13, 15, 14, 14, 14, 13, 13, 13, 14, 18, 18, 21, 19, 22, 21, 21, 22, 24, 22, 24, 24, 28, 28, 28, 27, 28, 26, 27, 27, 26, 25, 27, 28, 33, 39, 45, 51, 53, 54, 57, 57, 45, 14, 21, 20, 19, 22, 17, 18, 19, 18, 58, 111, 112, 110, 113, 109, 111, 112, 112, 110,
		110, 109, 111, 107, 110, 106, 110, 109, 109, 107, 109, 109, 109, 108, 111, 109, 111, 111, 109, 110, 112, 112, 112, 109, 113, 108, 111, 108, 112, 110, 144, 178, 167, 168, 173, 169, 172, 173, 173, 173, 173, 170, 174, 173, 176, 182, 195, 190, 189, 189, 121, 97, 120, 168, 172, 167, 168, 201, 192, 192, 187, 185, 170, 171, 188, 160, 181, 158, 192, 177, 192, 198, 206, 198, 192, 194, 145, 96, 147, 183, 92, 127, 189, 135, 115, 145, 186, 168, 178, 173, 127, 72, 116, 156, 184, 170, 173, 175, 171, 130, 94, 113, 106, 107, 107, 106, 106, 103, 106, 104, 105, 102, 103, 103, 101, 100, 100, 97, 99, 98, 99, 97, 96, 94, 96, 96, 93, 42, 37, 37, 18, 7, 14, 10, 11, 10, 11, 12, 12, 12, 12, 11, 14, 14, 18, 17, 17, 15, 18, 17, 19, 16, 16, 12, 15, 12, 13, 10, 12, 19, 43, 72, 63, 41, 35, 33, 35, 35, 34, 32, 34, 32, 35, 32, 34, 32, 33, 33, 33, 32, 34, 32, 34, 32, 36, 50, 74, 84, 88, 89, 91, 88, 85, 77, 68, 53, 45, 37, 35, 31, 32, 28, 30, 28, 31, 30, 30, 27, 27, 19, 12, 11, 9, 7, 9, 9, 9, 9, 12, 30, 54, 59, 75, 67, 73, 66, 69, 67, 69, 67, 68, 68, 70, 68, 71, 69, 68, 69, 72, 67, 66, 58, 41, 58, 51, 45, 50, 69, 73, 69, 70, 71, 75, 74, 76, 76, 76, 75, 75, 73, 78, 78, 79, 77, 75, 77, 77, 75, 77, 76, 67, 46, 47, 47, 48, 46, 48, 45, 48, 46, 48, 46, 47, 46, 47, 46, 47, 45, 48, 46, 47, 45, 47, 48, 55, 57, 60, 59, 61, 60, 59, 58, 59, 57, 60, 58, 60, 58, 58, 56, 59, 56, 57, 54, 55, 53, 52, 50, 48, 24,
		23, 15, 12, 14, 14, 13, 14, 13, 13, 12, 13, 13, 18, 20, 21, 20, 23, 22, 22, 21, 23, 21, 23, 23, 24, 25, 29, 31, 32, 30, 33, 32, 34, 33, 37, 40, 48, 52, 58, 57, 53, 43, 40, 50, 45, 17, 13, 20, 26, 23, 16, 17, 19, 17, 55, 110, 111, 111, 113, 110, 113, 114, 113, 112, 111, 111, 112, 108, 109, 107, 108, 110, 110, 109, 111, 109, 109, 109, 111, 108, 109, 111, 110, 109, 112, 110, 112, 111, 110, 110, 109, 107, 111, 110, 138, 178, 167, 169, 173, 169, 173, 172, 173, 171, 172, 173, 172, 175, 176, 182, 192, 190, 191, 188, 123, 129, 105, 162, 182, 150, 169, 197, 185, 183, 173, 194, 187, 189, 188, 172, 173, 173, 193, 181, 188, 202, 206, 202, 194, 191, 193, 187, 189, 190, 190, 190, 195, 147, 101, 149, 185, 167, 178, 173, 159, 105, 116, 181, 175, 173, 175, 173, 172, 131, 97, 112, 107, 106, 108, 106, 107, 103, 107, 104, 105, 102, 103, 102, 102, 99, 97, 97, 99, 97, 98, 96, 96, 96, 95, 95, 90, 43, 38, 37, 18, 5, 14, 13, 12, 12, 11, 10, 12, 10, 12, 9, 13, 13, 17, 22, 14, 15, 14, 14, 15, 14, 17, 15, 19, 20, 16, 10, 12, 19, 44, 74, 62, 40, 37, 34, 34, 33, 33, 31, 36, 33, 33, 33, 34, 33, 34, 33, 35, 32, 33, 31, 33, 32, 35, 50, 73, 82, 89, 88, 90, 86, 79, 69, 56, 45, 39, 32, 33, 29, 30, 29, 28, 29, 28, 28, 31, 27, 27, 19, 13, 10, 10, 7, 9, 7, 9, 8, 14, 32, 53, 56, 77, 68, 72, 69, 69, 70, 68, 67, 67, 69, 69, 69, 71, 69, 69, 71, 69, 67, 66, 58, 42, 59, 52, 44, 49, 70, 73, 69, 72, 71, 75, 73, 77, 76,
		21, 14, 13, 13, 13, 13, 13, 13, 13, 12, 13, 14, 15, 16, 17, 19, 19, 20, 20, 22, 40, 62, 79, 88, 94, 99, 103, 107, 110, 112, 117, 122, 122, 104, 96, 189, 112, 33, 24, 16, 14, 16, 17, 17, 17, 55, 108, 112, 111, 111, 111, 112, 113, 112, 111, 110, 110, 109, 108, 108, 110, 110, 109, 111, 108, 109, 109, 109, 109, 109, 109, 109, 111, 110, 109, 111, 108, 108, 124, 172, 167, 169, 172, 173, 172, 173, 172, 173, 173, 173, 177, 189, 194, 192, 190, 149, 125, 152, 181, 159, 172, 192, 182, 183, 194, 183, 191, 175, 164, 161, 192, 190, 191, 200, 202, 196, 195, 193, 193, 189, 189, 190, 190, 190, 188, 174, 175, 176, 141, 110, 119, 169, 178, 174, 175, 163, 116, 104, 108, 107, 107, 106, 107, 107, 106, 106, 104, 103, 102, 102, 100, 99, 97, 97, 96, 97, 96, 96, 95, 54, 36, 32, 13, 10, 11, 11, 10, 10, 10, 9, 11, 11, 10, 12, 12, 12, 11, 13, 16, 17, 20, 25, 23, 17, 15, 35, 37, 57, 66, 42, 35, 33, 34, 33, 33, 34, 33, 34, 33, 32, 34, 33, 34, 33, 32, 32, 34, 45, 66, 78, 78, 66, 54, 45, 37, 33, 31, 30, 30, 29, 30, 28, 28, 28, 27, 28, 26, 23, 15, 10, 9, 8, 8, 9, 8, 14, 33, 55, 69, 69, 70, 69, 70, 69, 65, 68, 69, 69, 71, 70, 70, 70, 70, 68, 58, 48, 58, 48, 50, 67, 72, 71, 71, 72, 73, 77, 77, 78, 75, 74, 77, 77, 78, 77, 77, 76, 76, 77, 69, 47, 47, 46, 46, 47, 46, 46, 46, 47, 47, 47, 47, 47, 47, 48, 45, 46, 46, 45, 46, 46, 47, 46, 46, 46, 44, 43, 43, 43, 43, 43, 45, 45, 45, 45, 45, 46, 45, 46, 45, 26,
		22, 15, 14, 14, 13, 13, 13, 13, 13, 11, 12, 10, 11, 12, 11, 13, 12, 13, 14, 13, 18, 25, 34, 39, 43, 47, 49, 52, 54, 56, 60, 66, 68, 68, 66, 137, 120, 31, 25, 21, 15, 15, 16, 16, 18, 53, 106, 110, 112, 111, 112, 111, 113, 113, 110, 112, 110, 108, 108, 106, 109, 110, 110, 111, 110, 109, 108, 109, 110, 108, 109, 109, 109, 108, 110, 111, 108, 108, 122, 171, 169, 172, 173, 173, 173, 174, 174, 174, 174, 174, 177, 188, 193, 191, 190, 180, 162, 176, 184, 170, 181, 190, 183, 180, 196, 189, 189, 180, 161, 170, 194, 193, 193, 201, 202, 196, 196, 195, 194, 190, 190, 190, 190, 190, 188, 174, 174, 175, 139, 140, 133, 166, 180, 172, 176, 163, 116, 106, 109, 107, 108, 105, 105, 107, 106, 106, 104, 103, 103, 103, 101, 99, 98, 97, 97, 98, 97, 96, 95, 56, 36, 34, 15, 11, 10, 10, 10, 10, 11, 10, 11, 11, 11, 13, 11, 11, 11, 13, 18, 21, 19, 22, 21, 21, 29, 43, 37, 58, 66, 42, 34, 34, 33, 33, 32, 34, 34, 34, 32, 31, 34, 33, 33, 33, 32, 34, 35, 46, 63, 69, 63, 52, 43, 37, 34, 33, 31, 31, 30, 30, 29, 28, 29, 28, 27, 27, 25, 22, 14, 10, 9, 8, 8, 8, 8, 15, 31, 56, 69, 69, 71, 70, 70, 69, 66, 68, 70, 70, 70, 70, 70, 70, 70, 68, 59, 48, 58, 49, 51, 68, 72, 72, 71, 72, 73, 76, 77, 78, 76, 74, 76, 77, 77, 76, 77, 77, 74, 77, 69, 48, 47, 47, 46, 46, 46, 46, 45, 47, 47, 46, 48, 46, 47, 47, 46, 46, 45, 46, 47, 47, 47, 46, 46, 45, 45, 46, 45, 44, 46, 46, 48, 46, 47, 47, 46, 47, 47, 48, 46, 27,
		23, 20, 17, 17, 15, 13, 13, 12, 13, 11, 11, 10, 11, 11, 10, 11, 10, 10, 10, 10, 11, 11, 13, 15, 17, 21, 20, 21, 22, 22, 23, 23, 24, 25, 23, 34, 33, 20, 21, 22, 21, 15, 16, 16, 16, 48, 103, 111, 113, 112, 112, 112, 111, 111, 110, 110, 108, 108, 110, 109, 107, 109, 111, 112, 110, 110, 110, 109, 110, 108, 110, 110, 109, 109, 109, 111, 109, 109, 120, 168, 173, 175, 175, 175, 172, 173, 172, 174, 175, 173, 179, 187, 192, 192, 191, 189, 175, 157, 188, 184, 187, 188, 183, 173, 195, 197, 189, 177, 162, 156, 190, 194, 191, 198, 202, 195, 195, 195, 196, 192, 189, 189, 191, 191, 189, 175, 172, 174, 134, 116, 124, 165, 180, 172, 176, 163, 116, 105, 108, 105, 109, 106, 107, 108, 107, 107, 105, 104, 104, 104, 101, 100, 98, 98, 96, 98, 97, 96, 94, 61, 34, 36, 19, 11, 9, 11, 12, 11, 10, 11, 12, 11, 11, 13, 12, 13, 10, 12, 18, 32, 30, 30, 31, 36, 42, 44, 36, 58, 67, 44, 34, 34, 34, 33, 33, 34, 33, 34, 32, 31, 34, 33, 33, 33, 32, 35, 35, 43, 55, 56, 51, 42, 36, 34, 33, 32, 30, 30, 31, 30, 31, 29, 28, 29, 27, 28, 25, 22, 14, 10, 9, 8, 9, 9, 8, 14, 28, 53, 70, 70, 71, 70, 70, 69, 67, 69, 69, 70, 70, 69, 70, 71, 71, 68, 60, 49, 56, 49, 51, 67, 74, 72, 72, 74, 73, 75, 77, 78, 76, 74, 76, 79, 78, 76, 78, 77, 76, 77, 69, 48, 47, 46, 47, 47, 45, 47, 46, 46, 46, 46, 47, 45, 46, 47, 46, 48, 47, 46, 47, 46, 48, 46, 46, 46, 47, 46, 45, 45, 46, 47, 47, 46, 46, 47, 48, 47, 47, 48, 47, 27,
		23, 26, 23, 22, 18, 13, 13, 13, 13, 11, 11, 10, 10, 10, 10, 11, 10, 10, 10, 9, 11, 10, 11, 11, 14, 15, 16, 17, 19, 18, 20, 18, 18, 19, 18, 20, 19, 18, 18, 20, 25, 19, 16, 17, 16, 45, 103, 111, 113, 113, 114, 112, 111, 111, 110, 110, 108, 108, 110, 108, 109, 108, 110, 111, 109, 111, 111, 111, 111, 110, 110, 109, 111, 111, 110, 111, 109, 110, 117, 167, 173, 174, 175, 175, 173, 175, 173, 173, 175, 175, 178, 187, 191, 191, 192, 155, 107, 149, 189, 188, 189, 191, 195, 187, 190, 189, 190, 177, 176, 173, 188, 195, 191, 196, 201, 195, 192, 193, 194, 194, 191, 189, 190, 191, 189, 177, 172, 174, 147, 102, 151, 176, 177, 175, 175, 164, 114, 105, 109, 106, 108, 108, 107, 107, 106, 106, 105, 104, 105, 104, 103, 101, 101, 99, 97, 98, 95, 96, 96, 60, 35, 36, 19, 11, 10, 11, 13, 12, 11, 11, 14, 12, 13, 13, 13, 11, 11, 13, 27, 47, 46, 46, 46, 47, 45, 43, 37, 59, 69, 45, 36, 34, 34, 35, 33, 34, 33, 32, 34, 33, 34, 34, 34, 34, 33, 34, 34, 37, 41, 43, 40, 35, 32, 31, 31, 32, 31, 30, 30, 29, 29, 28, 28, 29, 28, 28, 25, 22, 15, 10, 9, 7, 8, 8, 7, 12, 23, 48, 69, 70, 71, 69, 69, 70, 68, 70, 69, 70, 71, 67, 70, 70, 71, 68, 60, 50, 56, 49, 49, 68, 73, 73, 74, 75, 74, 74, 77, 77, 76, 74, 77, 78, 78, 77, 77, 77, 77, 77, 69, 47, 47, 47, 46, 46, 46, 46, 45, 46, 47, 46, 47, 45, 45, 46, 46, 47, 46, 47, 47, 46, 49, 47, 48, 48, 45, 47, 46, 46, 46, 45, 47, 45, 45, 47, 46, 48, 48, 48, 48, 28,
		22, 26, 24, 21, 19, 13, 13, 13, 13, 11, 11, 10, 10, 11, 10, 10, 10, 10, 9, 9, 10, 10, 10, 11, 12, 13, 12, 14, 16, 17, 19, 18, 19, 18, 18, 19, 19, 18, 18, 17, 22, 23, 20, 17, 15, 41, 101, 113, 114, 112, 115, 113, 113, 112, 109, 109, 108, 108, 108, 107, 109, 109, 109, 110, 109, 111, 108, 108, 112, 110, 108, 108, 110, 110, 109, 111, 110, 109, 115, 162, 174, 174, 175, 176, 175, 175, 174, 174, 175, 175, 179, 187, 192, 191, 191, 175, 148, 147, 187, 185, 193, 193, 199, 198, 193, 189, 189, 174, 166, 162, 190, 195, 201, 194, 202, 192, 191, 194, 194, 193, 190, 190, 190, 190, 188, 178, 174, 175, 130, 112, 117, 173, 178, 174, 177, 163, 114, 105, 109, 107, 108, 108, 107, 108, 105, 106, 106, 106, 104, 103, 103, 100, 99, 99, 98, 98, 96, 96, 95, 60, 35, 35, 17, 11, 10, 12, 12, 11, 11, 13, 14, 14, 16, 15, 14, 13, 12, 22, 41, 48, 50, 49, 48, 48, 46, 43, 38, 58, 67, 43, 35, 34, 34, 35, 33, 34, 32, 32, 33, 33, 33, 33, 33, 34, 33, 33, 32, 34, 36, 36, 35, 34, 32, 31, 31, 33, 31, 30, 31, 29, 29, 28, 28, 28, 27, 28, 25, 22, 14, 11, 10, 8, 9, 9, 8, 12, 21, 45, 68, 70, 71, 69, 70, 69, 66, 68, 69, 69, 70, 67, 69, 69, 70, 67, 61, 50, 57, 49, 48, 70, 72, 72, 74, 74, 74, 76, 77, 77, 76, 72, 74, 76, 77, 77, 77, 76, 77, 76, 67, 46, 47, 47, 47, 46, 45, 47, 46, 47, 47, 47, 47, 45, 47, 46, 46, 48, 47, 48, 48, 47, 49, 47, 48, 48, 46, 47, 47, 47, 47, 45, 47, 45, 45, 46, 46, 47, 46, 47, 47, 27
	);
	
	constant buffer_right : t_array_image := (
		18, 6, 4, 6, 5, 5, 5, 6, 5, 6, 5, 5, 5, 6, 6, 6, 5, 5, 5, 6, 5, 5, 6, 5, 7, 6, 7, 6, 7, 6, 6, 6, 8, 9, 11, 11, 13, 14, 19, 27, 38, 35, 28, 23, 29, 43, 54, 54, 55, 55, 56, 55, 56, 57, 62, 66, 75, 65, 63, 65, 44, 39, 39, 56, 43, 0, 10, 9, 8, 7, 6, 6, 7, 7, 9, 9, 7, 7, 10, 14, 16, 16, 16, 15, 18, 18, 22, 22, 23, 23, 24, 23, 24, 23, 24, 25, 27, 27, 26, 27, 38, 60, 55, 56, 57, 55, 57, 56, 55, 55, 55, 54, 54, 51, 53, 53, 54, 55, 55, 53, 56, 56, 55, 55, 55, 55, 54, 53, 55, 54, 55, 54, 54, 54, 55, 55, 55, 55, 55, 66, 93, 82, 86, 84, 86, 86, 87, 85, 86, 84, 85, 86, 86, 85, 89, 94, 95, 95, 95, 55, 35, 54, 93, 86, 76, 81, 100, 92, 80, 84, 97, 78, 93, 83, 90, 73, 89, 91, 90, 99, 105, 94, 99, 96, 97, 63, 53, 73, 98, 49, 61, 101, 77, 52, 64, 91, 86, 89, 86, 74, 56, 66, 78, 90, 84, 86, 87, 86, 69, 46, 55, 52, 51, 53, 54, 51, 52, 51, 50, 51, 50, 51, 51, 49, 51, 48, 49, 48, 48, 48, 48, 48, 47, 47, 48, 43, 20, 18, 13, 4, 5, 5, 10, 19, 37, 34, 23, 18, 17, 16, 16, 16, 17, 14, 16, 16, 17, 15, 17, 15, 17, 15, 16, 15, 15, 15, 17, 17, 22, 33, 42, 44, 45, 43, 42, 43, 43, 41, 40, 38, 36, 32, 26, 22, 20, 16, 15, 14, 15, 14, 14, 12, 12, 7, 6, 4, 4, 4, 4, 3, 4, 3, 4, 4, 5, 4, 6, 5, 5, 7, 13, 22, 29, 31, 35, 34, 35, 34, 33, 33,
		34, 31, 33, 34, 35, 34, 35, 33, 34, 33, 35, 33, 31, 28, 13, 6, 9, 8, 20, 29, 26, 24, 23, 26, 35, 35, 35, 35, 36, 35, 36, 38, 38, 37, 37, 37, 38, 37, 38, 37, 38, 37, 39, 37, 39, 37, 38, 33, 25, 22, 23, 22, 21, 22, 21, 21, 22, 22, 23, 23, 31, 38, 43, 22, 32, 14, 10, 11, 12, 11, 12, 11, 11, 11, 11, 11, 12, 11, 12, 11, 12, 11, 12, 12, 13, 12, 13, 12, 14, 13, 15, 14, 14, 13, 14, 14, 17, 20, 23, 22, 26, 25, 27, 38, 51, 56, 47, 40, 59, 85, 100, 100, 101, 99, 103, 99, 99, 102, 116, 126, 167, 156, 108, 155, 93, 17, 41, 48, 42, 16, 18, 24, 22, 13, 16, 12, 16, 15, 19, 18, 17, 14, 27, 44, 46, 45, 47, 45, 49, 49, 50, 49, 50, 49, 50, 51, 49, 48, 50, 49, 56, 57, 55, 53, 77, 122, 113, 114, 114, 110, 115, 115, 113, 112, 113, 110, 109, 108, 109, 110, 112, 108, 112, 110, 111, 111, 112, 109, 109, 109, 110, 110, 112, 111, 110, 110, 110, 109, 111, 111, 110, 111, 111, 134, 184, 169, 175, 170, 174, 172, 173, 174, 173, 171, 172, 173, 174, 175, 183, 190, 190, 190, 191, 138, 114, 130, 191, 173, 155, 170, 200, 184, 163, 175, 191, 159, 172, 183, 188, 163, 173, 187, 178, 196, 205, 198, 193, 196, 197, 131, 110, 194, 180, 99, 122, 198, 150, 92, 125, 186, 170, 178, 174, 139, 91, 127, 155, 186, 171, 174, 175, 170, 136, 95, 110, 103, 105, 105, 108, 104, 106, 105, 104, 103, 104, 102, 104, 101, 101, 96, 97, 97, 98, 98, 95, 95, 95, 95, 96, 89, 42, 36, 24, 9, 12, 11, 23, 42, 75, 67, 47, 36, 37, 34, 35, 33, 33, 32, 34, 33,
		34, 32, 33, 32, 32, 32, 33, 30, 33, 33, 32, 34, 45, 66, 84, 88, 90, 86, 86, 84, 85, 83, 80, 74, 70, 56, 48, 40, 36, 31, 31, 27, 29, 29, 27, 25, 22, 14, 12, 8, 8, 8, 10, 8, 10, 8, 10, 8, 10, 10, 13, 12, 14, 13, 27, 45, 55, 62, 73, 68, 70, 69, 69, 69, 66, 63, 69, 68, 69, 69, 69, 68, 69, 68, 72, 67, 65, 57, 24, 12, 17, 17, 43, 59, 54, 48, 46, 54, 73, 70, 74, 68, 71, 71, 71, 76, 77, 74, 75, 74, 76, 75, 78, 76, 77, 74, 80, 76, 77, 75, 75, 66, 51, 45, 45, 46, 44, 44, 44, 44, 44, 43, 45, 48, 60, 75, 80, 41, 27, 13, 8, 12, 12, 11, 13, 11, 12, 11, 11, 12, 13, 11, 13, 11, 12, 11, 11, 12, 12, 11, 14, 12, 14, 12, 14, 13, 15, 13, 14, 14, 18, 19, 22, 21, 22, 21, 25, 25, 29, 31, 34, 34, 45, 60, 66, 64, 64, 62, 64, 60, 57, 56, 68, 81, 106, 142, 61, 109, 74, 14, 44, 51, 42, 17, 23, 37, 24, 14, 16, 14, 16, 15, 17, 17, 17, 14, 26, 51, 47, 49, 50, 48, 50, 48, 50, 49, 50, 50, 51, 48, 50, 47, 51, 50, 54, 57, 58, 52, 77, 117, 113, 116, 115, 110, 113, 113, 114, 111, 111, 109, 108, 107, 108, 110, 112, 109, 111, 112, 112, 110, 111, 107, 108, 107, 112, 108, 112, 111, 111, 110, 111, 109, 109, 108, 108, 109, 111, 129, 183, 169, 173, 171, 173, 172, 173, 173, 174, 171, 173, 170, 173, 175, 182, 190, 192, 191, 193, 175, 119, 131, 164, 196, 140, 179, 201, 187, 165, 175, 194, 175, 191, 191, 173, 155, 172, 188, 178, 194, 199, 207, 194, 190, 198, 150, 72, 151, 193, 96, 122, 200,
		146, 88, 119, 186, 170, 178, 173, 122, 86, 121, 140, 195, 165, 176, 175, 171, 136, 95, 109, 103, 106, 105, 106, 103, 107, 106, 107, 103, 106, 103, 104, 103, 102, 98, 99, 96, 99, 96, 98, 94, 96, 95, 97, 89, 39, 37, 24, 9, 11, 10, 22, 43, 73, 69, 45, 37, 35, 34, 36, 32, 33, 33, 34, 33, 33, 32, 34, 31, 32, 32, 32, 32, 34, 32, 33, 31, 47, 67, 85, 88, 89, 87, 86, 82, 87, 85, 77, 65, 56, 46, 40, 34, 31, 30, 30, 29, 28, 30, 29, 26, 22, 13, 12, 8, 9, 8, 9, 7, 9, 8, 9, 8, 10, 10, 13, 12, 14, 14, 25, 44, 57, 65, 72, 69, 71, 68, 70, 69, 69, 66, 68, 68, 71, 68, 68, 67, 70, 71, 72, 67, 66, 57, 24, 10, 15, 17, 46, 60, 52, 47, 43, 55, 72, 71, 71, 70, 72, 71, 74, 75, 76, 74, 77, 75, 75, 75, 77, 76, 77, 75, 78, 75, 75, 73, 75, 66, 50, 45, 47, 45, 46, 41, 45, 45, 46, 45, 46, 48, 59, 66, 70, 35, 26, 13, 10, 12, 12, 11, 12, 11, 12, 11, 11, 11, 12, 11, 11, 11, 12, 11, 13, 11, 13, 12, 12, 12, 15, 12, 14, 13, 14, 12, 14, 13, 16, 18, 23, 20, 22, 23, 23, 22, 26, 27, 28, 30, 36, 46, 47, 44, 41, 38, 37, 35, 33, 31, 30, 31, 35, 37, 40, 41, 44, 43, 51, 55, 48, 17, 21, 51, 37, 12, 14, 15, 14, 16, 17, 17, 18, 15, 21, 51, 49, 48, 49, 49, 50, 48, 50, 51, 52, 50, 52, 50, 51, 49, 51, 51, 56, 58, 60, 52, 69, 117, 110, 114, 114, 112, 114, 112, 112, 109, 110, 107, 108, 107, 110, 109, 111, 110, 110, 111, 112, 110, 110, 108, 110, 108, 111, 108,
		110, 109, 111, 110, 109, 109, 109, 109, 108, 106, 111, 125, 181, 170, 172, 169, 172, 172, 173, 172, 173, 171, 174, 173, 175, 174, 180, 190, 191, 190, 189, 145, 84, 108, 174, 190, 152, 164, 205, 187, 171, 169, 201, 177, 157, 187, 172, 157, 168, 190, 176, 193, 199, 209, 200, 188, 195, 165, 146, 170, 194, 148, 114, 204, 159, 108, 140, 183, 169, 177, 174, 128, 109, 94, 148, 186, 171, 172, 174, 173, 137, 93, 112, 104, 105, 104, 105, 105, 105, 104, 107, 104, 105, 104, 102, 103, 103, 97, 99, 97, 100, 99, 96, 96, 97, 96, 98, 89, 43, 38, 26, 8, 12, 11, 22, 40, 71, 69, 47, 36, 34, 35, 36, 34, 34, 32, 34, 33, 36, 32, 33, 34, 34, 34, 34, 33, 34, 33, 34, 33, 46, 66, 83, 88, 89, 88, 87, 86, 86, 81, 70, 55, 47, 39, 34, 30, 30, 30, 30, 29, 29, 28, 29, 26, 23, 13, 11, 8, 9, 9, 8, 8, 9, 7, 9, 9, 8, 11, 13, 12, 15, 14, 25, 40, 56, 63, 73, 68, 70, 68, 69, 69, 70, 67, 68, 68, 70, 68, 69, 68, 69, 69, 72, 67, 67, 56, 25, 9, 15, 18, 44, 59, 52, 44, 44, 53, 70, 69, 71, 68, 71, 71, 75, 76, 77, 74, 76, 74, 76, 75, 77, 76, 77, 73, 77, 75, 76, 76, 76, 67, 51, 45, 46, 46, 46, 44, 46, 44, 47, 44, 47, 46, 52, 55, 59, 30, 23, 14, 10, 12, 12, 11, 12, 12, 11, 12, 11, 10, 13, 10, 11, 9, 12, 10, 12, 11, 13, 12, 14, 13, 16, 13, 14, 12, 14, 13, 14, 13, 17, 19, 20, 20, 22, 21, 22, 23, 24, 24, 25, 25, 28, 32, 33, 29, 30, 29, 28, 27, 27, 26, 28, 26, 30, 33, 38, 44, 51, 54, 56, 57,
		48, 14, 25, 16, 24, 21, 15, 13, 15, 16, 16, 16, 18, 16, 18, 49, 52, 50, 49, 49, 50, 48, 50, 50, 50, 53, 55, 53, 54, 50, 50, 52, 57, 59, 60, 54, 67, 112, 113, 112, 112, 111, 112, 111, 111, 109, 110, 109, 109, 107, 110, 108, 110, 107, 109, 107, 109, 108, 109, 109, 111, 111, 111, 108, 110, 107, 109, 109, 110, 110, 110, 109, 110, 108, 110, 122, 181, 172, 173, 170, 174, 172, 175, 173, 174, 171, 173, 172, 176, 174, 180, 192, 193, 187, 189, 168, 95, 120, 180, 184, 154, 173, 198, 195, 181, 177, 195, 159, 160, 182, 172, 185, 172, 178, 188, 187, 200, 206, 204, 190, 196, 158, 92, 131, 196, 98, 112, 181, 145, 137, 169, 178, 171, 177, 175, 139, 95, 120, 157, 185, 171, 173, 176, 172, 134, 94, 111, 106, 105, 106, 106, 103, 103, 103, 105, 102, 103, 103, 103, 102, 101, 98, 98, 97, 100, 98, 98, 94, 96, 95, 97, 90, 44, 37, 25, 9, 12, 11, 22, 39, 68, 69, 46, 36, 36, 33, 36, 34, 34, 33, 34, 34, 33, 33, 35, 33, 34, 32, 34, 33, 34, 33, 32, 33, 43, 64, 82, 86, 88, 88, 90, 85, 81, 72, 60, 45, 39, 34, 33, 31, 29, 28, 29, 28, 30, 29, 29, 27, 23, 14, 11, 9, 8, 9, 9, 9, 9, 8, 9, 8, 10, 10, 14, 13, 13, 14, 22, 40, 54, 59, 75, 68, 70, 69, 70, 67, 69, 68, 68, 67, 71, 68, 70, 68, 69, 69, 70, 66, 65, 58, 25, 9, 17, 19, 43, 58, 51, 45, 45, 52, 71, 70, 71, 69, 73, 72, 74, 75, 75, 75, 75, 73, 74, 75, 79, 77, 78, 74, 76, 75, 75, 75, 78, 66, 52, 43, 46, 45, 47, 43, 45, 45, 47, 44, 47, 45, 48, 50, 52, 26,
		22, 14, 10, 11, 12, 11, 11, 12, 12, 12, 13, 11, 12, 11, 11, 11, 12, 11, 12, 11, 13, 12, 14, 12, 14, 12, 14, 13, 13, 12, 13, 12, 15, 19, 23, 21, 22, 19, 23, 21, 24, 22, 22, 23, 26, 24, 29, 27, 29, 27, 29, 26, 27, 25, 30, 30, 36, 41, 49, 53, 56, 53, 54, 55, 46, 14, 17, 21, 25, 25, 19, 13, 15, 14, 16, 16, 20, 17, 16, 37, 58, 47, 52, 51, 50, 51, 51, 49, 49, 50, 53, 52, 53, 51, 52, 54, 61, 61, 63, 54, 66, 113, 113, 113, 115, 110, 112, 113, 112, 111, 110, 109, 110, 106, 108, 107, 109, 109, 110, 106, 110, 107, 108, 108, 109, 108, 111, 110, 111, 109, 114, 111, 112, 110, 112, 109, 108, 109, 111, 120, 174, 172, 170, 172, 172, 171, 174, 172, 173, 172, 174, 173, 176, 176, 183, 192, 193, 190, 193, 136, 131, 138, 129, 194, 155, 172, 190, 189, 194, 174, 197, 186, 189, 187, 173, 165, 170, 195, 185, 185, 201, 204, 204, 191, 193, 180, 169, 175, 193, 170, 177, 192, 161, 97, 151, 183, 171, 176, 174, 149, 85, 128, 176, 174, 173, 174, 175, 173, 133, 96, 112, 104, 105, 106, 106, 103, 104, 105, 104, 103, 102, 101, 101, 100, 99, 96, 97, 96, 97, 98, 98, 94, 97, 94, 96, 87, 43, 38, 29, 11, 12, 13, 24, 39, 71, 67, 46, 38, 36, 35, 34, 34, 35, 33, 34, 33, 34, 34, 34, 33, 34, 33, 34, 32, 34, 33, 33, 34, 44, 65, 81, 86, 88, 88, 89, 81, 73, 60, 49, 38, 34, 32, 31, 29, 29, 28, 28, 27, 30, 31, 29, 25, 22, 13, 12, 8, 9, 7, 9, 8, 10, 7, 9, 8, 11, 10, 13, 12, 14, 13, 21, 41, 52, 57, 73, 67, 71, 68, 70, 68,
		21, 12, 10, 12, 11, 12, 12, 11, 11, 11, 12, 11, 11, 12, 12, 12, 12, 12, 13, 12, 13, 13, 13, 13, 12, 13, 12, 15, 18, 19, 23, 23, 23, 24, 24, 26, 32, 54, 80, 97, 107, 112, 118, 124, 128, 134, 136, 142, 146, 144, 95, 107, 129, 56, 25, 15, 13, 17, 21, 18, 19, 18, 16, 16, 17, 17, 20, 47, 58, 56, 56, 56, 56, 57, 56, 57, 57, 59, 59, 59, 62, 60, 58, 58, 99, 114, 113, 113, 113, 113, 113, 111, 111, 110, 109, 109, 109, 109, 109, 108, 109, 108, 108, 109, 109, 109, 109, 109, 110, 108, 111, 109, 109, 109, 107, 110, 132, 171, 171, 169, 175, 173, 174, 173, 173, 175, 174, 175, 180, 191, 194, 193, 177, 121, 133, 145, 186, 157, 184, 186, 179, 185, 192, 192, 190, 168, 168, 175, 193, 184, 198, 201, 199, 196, 193, 193, 191, 189, 189, 191, 190, 190, 181, 175, 174, 167, 119, 106, 139, 181, 171, 175, 173, 142, 101, 109, 106, 106, 105, 106, 107, 104, 104, 103, 101, 102, 100, 100, 100, 96, 96, 95, 96, 96, 95, 95, 74, 39, 32, 14, 37, 41, 36, 60, 69, 41, 36, 34, 34, 32, 33, 33, 34, 34, 33, 34, 34, 34, 33, 33, 33, 33, 34, 43, 64, 78, 77, 67, 55, 45, 37, 33, 31, 29, 29, 30, 29, 29, 29, 28, 27, 28, 26, 23, 15, 10, 8, 8, 9, 7, 9, 8, 9, 9, 10, 13, 13, 14, 16, 30, 53, 65, 71, 69, 68, 69, 69, 67, 66, 69, 69, 69, 70, 69, 69, 71, 68, 63, 36, 13, 17, 29, 54, 55, 48, 47, 61, 71, 70, 70, 71, 72, 75, 76, 77, 76, 73, 75, 76, 76, 76, 75, 76, 75, 75, 75, 60, 47, 46, 46, 47, 46, 46, 46, 46, 46, 45, 45, 46, 26,
		21, 13, 11, 12, 11, 11, 11, 11, 11, 11, 12, 12, 12, 12, 11, 12, 12, 13, 13, 12, 13, 13, 13, 13, 12, 13, 11, 12, 12, 13, 15, 15, 15, 16, 15, 17, 20, 33, 53, 69, 79, 83, 89, 94, 97, 100, 104, 113, 120, 122, 120, 169, 219, 118, 26, 27, 14, 14, 20, 19, 21, 21, 16, 17, 16, 19, 18, 38, 59, 58, 57, 57, 57, 57, 57, 59, 58, 60, 61, 60, 60, 59, 58, 58, 99, 115, 112, 112, 112, 112, 113, 113, 111, 111, 109, 109, 108, 108, 110, 110, 111, 110, 110, 109, 109, 110, 109, 109, 109, 107, 111, 109, 109, 110, 108, 109, 130, 170, 171, 170, 176, 173, 174, 174, 174, 176, 174, 175, 181, 192, 194, 193, 187, 158, 146, 174, 178, 162, 184, 188, 179, 185, 194, 189, 191, 165, 158, 179, 195, 190, 199, 202, 200, 196, 194, 194, 192, 190, 189, 189, 191, 189, 182, 173, 175, 168, 125, 124, 146, 179, 175, 173, 174, 141, 103, 110, 106, 106, 106, 104, 106, 105, 104, 103, 102, 103, 102, 101, 100, 97, 97, 96, 96, 96, 96, 95, 77, 41, 33, 26, 45, 40, 35, 60, 69, 43, 36, 35, 34, 33, 34, 34, 33, 34, 33, 33, 34, 34, 33, 33, 33, 34, 36, 45, 61, 70, 64, 53, 44, 37, 34, 32, 30, 28, 29, 29, 29, 28, 28, 28, 28, 27, 26, 23, 15, 11, 9, 8, 9, 7, 9, 8, 9, 9, 10, 14, 13, 13, 16, 28, 54, 66, 70, 70, 69, 69, 69, 67, 66, 69, 70, 70, 69, 69, 69, 71, 68, 62, 35, 12, 17, 29, 53, 55, 47, 47, 62, 73, 72, 72, 72, 73, 75, 76, 76, 76, 74, 74, 77, 78, 76, 76, 77, 75, 75, 75, 60, 47, 46, 45, 47, 45, 46, 46, 45, 45, 45, 45, 46, 26,
		21, 12, 11, 12, 11, 12, 11, 11, 12, 11, 13, 11, 11, 12, 10, 12, 12, 13, 15, 13, 15, 13, 13, 13, 12, 12, 11, 11, 11, 10, 11, 10, 11, 11, 10, 12, 11, 13, 16, 19, 25, 28, 29, 31, 31, 32, 33, 36, 38, 39, 42, 52, 71, 45, 18, 26, 18, 14, 17, 19, 16, 18, 20, 22, 15, 19, 16, 27, 56, 55, 58, 58, 57, 58, 58, 59, 59, 60, 61, 59, 60, 60, 58, 60, 97, 114, 114, 113, 112, 112, 113, 112, 110, 110, 110, 107, 108, 108, 107, 109, 111, 111, 110, 108, 109, 111, 111, 109, 110, 109, 109, 109, 110, 111, 108, 110, 129, 172, 176, 174, 177, 173, 174, 174, 174, 176, 175, 176, 181, 191, 194, 194, 192, 190, 182, 179, 191, 185, 189, 188, 180, 181, 200, 193, 188, 173, 159, 174, 194, 192, 195, 203, 199, 197, 196, 195, 195, 190, 189, 191, 191, 189, 182, 173, 174, 163, 123, 137, 142, 183, 172, 173, 173, 138, 102, 110, 105, 105, 107, 104, 107, 105, 106, 104, 104, 103, 102, 102, 100, 99, 97, 96, 96, 96, 95, 95, 74, 41, 39, 42, 46, 40, 35, 61, 68, 43, 36, 34, 34, 33, 34, 33, 34, 34, 32, 32, 33, 34, 34, 33, 34, 34, 35, 43, 53, 56, 50, 43, 36, 33, 33, 32, 31, 30, 29, 29, 29, 30, 29, 28, 30, 27, 26, 23, 15, 11, 8, 9, 9, 9, 9, 8, 9, 10, 11, 13, 13, 13, 14, 24, 52, 66, 71, 70, 69, 69, 68, 68, 67, 68, 70, 70, 69, 69, 70, 70, 67, 62, 34, 13, 16, 30, 54, 54, 47, 47, 62, 73, 72, 72, 73, 72, 74, 76, 77, 76, 74, 75, 78, 78, 77, 77, 77, 76, 76, 75, 59, 46, 47, 46, 47, 45, 46, 46, 46, 47, 45, 46, 46, 27,
		22, 12, 10, 11, 10, 11, 11, 11, 11, 10, 12, 11, 11, 12, 11, 12, 13, 16, 21, 21, 19, 19, 14, 13, 12, 12, 11, 10, 10, 10, 10, 9, 10, 10, 9, 11, 10, 10, 10, 10, 14, 16, 17, 18, 17, 19, 19, 19, 19, 19, 20, 20, 19, 18, 16, 21, 23, 19, 15, 16, 18, 17, 26, 37, 15, 20, 17, 19, 46, 57, 59, 57, 57, 57, 57, 59, 59, 58, 59, 58, 59, 59, 57, 57, 95, 114, 114, 114, 114, 112, 111, 109, 110, 110, 107, 109, 111, 110, 107, 107, 110, 110, 110, 110, 110, 110, 109, 109, 110, 110, 111, 110, 110, 110, 109, 110, 126, 169, 176, 175, 178, 174, 175, 173, 172, 175, 174, 176, 181, 192, 193, 192, 188, 161, 115, 161, 199, 187, 191, 190, 190, 180, 193, 196, 186, 173, 171, 175, 192, 193, 191, 201, 200, 194, 194, 194, 194, 192, 190, 188, 191, 190, 183, 174, 173, 169, 119, 110, 165, 177, 176, 174, 174, 138, 100, 110, 105, 105, 107, 105, 106, 106, 105, 105, 103, 103, 103, 102, 100, 100, 98, 96, 97, 95, 95, 96, 77, 41, 43, 47, 46, 40, 36, 61, 70, 43, 35, 34, 34, 34, 33, 33, 34, 33, 33, 33, 33, 34, 34, 33, 33, 32, 34, 38, 41, 43, 40, 36, 34, 32, 31, 32, 32, 31, 29, 30, 29, 29, 29, 29, 28, 26, 25, 23, 14, 10, 9, 8, 8, 7, 9, 8, 8, 9, 10, 14, 14, 13, 14, 20, 47, 67, 72, 71, 70, 70, 69, 67, 68, 68, 69, 69, 68, 68, 69, 71, 68, 61, 33, 12, 18, 30, 54, 54, 46, 46, 62, 73, 72, 73, 73, 73, 73, 76, 77, 76, 75, 74, 76, 77, 76, 75, 77, 76, 77, 74, 59, 47, 47, 46, 46, 46, 46, 47, 46, 48, 46, 46, 46, 26,
		22, 12, 11, 12, 11, 11, 11, 11, 11, 11, 12, 11, 11, 12, 11, 12, 12, 15, 24, 25, 21, 21, 14, 13, 12, 13, 11, 10, 10, 9, 10, 9, 10, 9, 10, 10, 9, 10, 9, 9, 12, 13, 13, 16, 17, 20, 18, 19, 18, 17, 19, 19, 20, 19, 17, 18, 21, 22, 18, 15, 19, 18, 33, 45, 22, 16, 18, 17, 34, 61, 55, 56, 56, 56, 57, 58, 57, 57, 57, 58, 58, 58, 57, 56, 92, 114, 115, 114, 114, 113, 113, 111, 110, 110, 108, 109, 108, 108, 109, 108, 109, 110, 110, 110, 110, 111, 111, 110, 109, 108, 112, 111, 110, 110, 109, 110, 124, 168, 176, 176, 177, 177, 176, 176, 175, 176, 176, 178, 181, 192, 192, 192, 187, 151, 133, 158, 197, 189, 191, 196, 205, 199, 190, 191, 188, 165, 164, 171, 191, 198, 199, 196, 199, 192, 193, 194, 194, 192, 190, 189, 190, 189, 184, 174, 174, 163, 103, 108, 149, 180, 173, 175, 174, 138, 100, 110, 106, 106, 107, 105, 106, 105, 104, 104, 104, 104, 102, 101, 100, 99, 98, 97, 97, 95, 95, 95, 77, 41, 43, 47, 46, 40, 37, 59, 69, 43, 36, 35, 35, 34, 34, 33, 33, 33, 34, 33, 33, 34, 34, 33, 33, 33, 33, 35, 36, 36, 34, 33, 33, 31, 32, 31, 31, 31, 29, 29, 28, 29, 28, 28, 27, 27, 25, 24, 15, 11, 9, 8, 8, 7, 8, 8, 9, 9, 11, 15, 14, 13, 13, 17, 42, 65, 71, 70, 69, 69, 68, 67, 66, 68, 69, 69, 68, 67, 67, 71, 67, 62, 33, 12, 17, 30, 54, 54, 47, 46, 62, 73, 72, 73, 74, 73, 74, 77, 76, 76, 74, 72, 74, 75, 75, 75, 76, 75, 75, 73, 59, 47, 46, 47, 46, 47, 46, 47, 46, 47, 47, 48, 47, 27
	);	

    -- Definicion de el tipo arreglo para La transpferencia de los datos entre los
    -- bufferes.
    type ARRAY_ASSIGN is array(0 to D - 1) of std_logic_vector(DATA_W downto 0);

    -- Declaraci?n de los registros que van a contener los datos que se van a 
    -- transferir entre los bufferes.
    signal assign : ARRAY_ASSIGN := (others => (others => '0')); 

    -- Decraraci?n de los registros que se usan para hacer el control de el procesado.
    signal enable_counter : std_logic := '0';
    signal enable_write_l : std_logic := '0';
    signal enable_write_r : std_logic_vector(D - 1 downto 0) := (others => '0');
    signal process_wait   : std_logic_vector(D - 1 downto 0) := (others => '0');
    signal cost_out       : COSTES;
    signal x_column       : std_logic_vector(COOR_W downto 0);
    signal y_row          : std_logic_vector(COOR_W downto 0);
    signal vs             : std_logic;

begin
    enable_counter <= adv and process_wait(0);

    addr_generator_inst : addr_generator
    port map(
        clk        => clk,
        rst        => rst,
        adv        => enable_counter,
        vs         => vs,
        column     => x_column,
        row        => y_row,
        addr_left  => addr_left,
        addr_right => addr_right,
        addr_out   => addr_out
    );
    
    processor_buffer_for : for i in 0 to D - 1 generate
        processor_buffer_insta : processor_buffer
        port map(
            clk          => clk,
            rst          => rst,
            adv          => adv,
            wrena_l      => enable_write_l,
            wrena_r      => enable_write_r(i),
            left         => pixel_left,
            right        => assign(i),
            row          => y_row,
            cost         => cost_out(i),
            process_wait => process_wait(i)
        );
    end generate;
	
	pixel_left <=  std_logic_vector(to_unsigned(buffer_left(to_integer(unsigned(addr_left))), 8));
	pixel_right <= std_logic_vector(to_unsigned(buffer_right(to_integer(unsigned(addr_right))), 8));

    assign_process : process(pixel_left, pixel_right)
    begin
		        case(x_column) is
                    when b"000000000" =>
                        enable_write_l <= '1';
                        enable_write_r <= x"0000000000000001";
                        assign(0) <= pixel_right;
                    when b"000000001" =>
                        enable_write_l <= '1';
                        enable_write_r <= x"0000000000000003";
                        for i in 0 to 1 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000000010" =>
                        enable_write_l <= '1';
                        enable_write_r <= x"0000000000000007";
                        for i in 0 to 2 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000000011" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"000000000000000E";
                        for i in 1 to 3 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000000100" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"000000000000001C";
                        for i in 2 to 4 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000000101" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000000000038";
                        for i in 3 to 5 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000000110" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000000000070";
                        for i in 4 to 6 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000000111" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"00000000000000E0";
                        for i in 5 to 7 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000001000" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"00000000000001C0";
                        for i in 6 to 8 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000001001" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000000000380";
                        for i in 7 to 9 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000001010" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000000000700";
                        for i in 8 to 10 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000001011" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000000000E00";
                        for i in 9 to 11 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000001100" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000000001C00";
                        for i in 10 to 12 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000001101" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000000003800";
                        for i in 11 to 13 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000001110" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000000007000";
                        for i in 12 to 14 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000001111" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"000000000000E000";
                        for i in 13 to 15 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000010000" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"000000000001C000";
                        for i in 14 to 16 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000010001" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000000038000";
                        for i in 15 to 17 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000010010" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000000070000";
                        for i in 16 to 18 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000010011" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"00000000000E0000";
                        for i in 17 to 19 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000010100" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"00000000001C0000";
                        for i in 18 to 20 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000010101" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000000380000";
                        for i in 19 to 21 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000010110" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000000700000";
                        for i in 20 to 22 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000010111" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000000E00000";
                        for i in 21 to 23 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000011000" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000001C00000";
                        for i in 22 to 24 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000011001" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000003800000";
                        for i in 23 to 25 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000011010" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000007000000";
                        for i in 24 to 26 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000011011" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"000000000E000000";
                        for i in 25 to 27 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000011100" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"000000001C000000";
                        for i in 26 to 28 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000011101" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000038000000";
                        for i in 27 to 29 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000011110" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000070000000";
                        for i in 28 to 30 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000011111" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"00000000E0000000";
                        for i in 29 to 31 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000100000" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"00000001C0000000";
                        for i in 30 to 32 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000100001" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000380000000";
                        for i in 31 to 33 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000100010" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000700000000";
                        for i in 32 to 34 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000100011" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000E00000000";
                        for i in 33 to 35 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000100100" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000001C00000000";
                        for i in 34 to 36 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000100101" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000380000000";
                        for i in 35 to 37 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000100110" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000007000000000";
                        for i in 36 to 38 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000100111" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"000000E000000000";
                        for i in 37 to 39 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000101000" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"000001C000000000";
                        for i in 38 to 40 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000101001" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000038000000000";
                        for i in 39 to 41 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000101010" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000070000000000";
                        for i in 40 to 42 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000101011" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"00000E0000000000";
                        for i in 41 to 43 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000101100" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"00001C0000000000";
                        for i in 42 to 44 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000101101" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000380000000000";
                        for i in 43 to 45 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000101110" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000700000000000";
                        for i in 44 to 46 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000101111" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000E00000000000";
                        for i in 45 to 47 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000110000" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0001C00000000000";
                        for i in 46 to 48 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000110001" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0003800000000000";
                        for i in 47 to 49 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000110010" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0007000000000000";
                        for i in 48 to 50 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000110011" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"000E000000000000";
                        for i in 49 to 51 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000110100" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"001C000000000000";
                        for i in 50 to 52 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000110101" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0038000000000000";
                        for i in 51 to 53 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000110110" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0070000000000000";
                        for i in 52 to 54 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000110111" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"00E0000000000000";
                        for i in 53 to 55 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000111000" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"01C0000000000000";
                        for i in 54 to 56 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000111001" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0380000000000000";
                        for i in 55 to 57 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000111010" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0700000000000000";
                        for i in 56 to 58 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000111011" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0E00000000000000";
                        for i in 57 to 59 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000111100" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"1C00000000000000";
                        for i in 58 to 60 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000111101" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"3800000000000000";
                        for i in 59 to 61 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000111110" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"7000000000000000";
                        for i in 60 to 62 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"000111111" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"E000000000000000";
                        for i in 61 to 63 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"001000000" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"C000000000000000";
                        for i in 62 to 63 loop
                            assign(i) <= pixel_right;
                        end loop;
                    when b"001000001" =>
                        enable_write_l <= '0';
                        enable_write_r <= x"8000000000000000";
                        assign(63) <= pixel_right;
                    when others =>
                        enable_write_l <= '0';
                        enable_write_r <= x"0000000000000000";
                        for i in 0 to D - 1 loop
                            assign(i) <= (others => '0');
                        end loop;
                end case;
--                    if x_column =  b"000000000" then
--                        enable_write_l <= '1';
--                        enable_write_r <= x"0000000000000001";
--                        assign(0) <= pixel_right;
--                    elsif x_column = b"000000001" then
--                        enable_write_l <= '1';
--                        enable_write_r <= x"0000000000000003";
--                        for i in 0 to 1 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000000010" then
--                        enable_write_l <= '1';
--                        enable_write_r <= x"0000000000000007";
--                        for i in 0 to 2 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000000011" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"000000000000000E";
--                        for i in 1 to 3 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000000100" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"000000000000001C";
--                        for i in 2 to 4 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000000101" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000000000038";
--                        for i in 3 to 5 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000000110" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000000000070";
--                        for i in 4 to 6 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000000111" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"00000000000000E0";
--                        for i in 5 to 7 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000001000" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"00000000000001C0";
--                        for i in 6 to 8 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000001001" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000000000380";
--                        for i in 7 to 9 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000001010" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000000000700";
--                        for i in 8 to 10 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000001011" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000000000E00";
--                        for i in 9 to 11 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000001100" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000000001C00";
--                        for i in 10 to 12 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000001101" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000000003800";
--                        for i in 11 to 13 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000001110" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000000007000";
--                        for i in 12 to 14 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000001111" then 
--                        enable_write_l <= '0';
--                        enable_write_r <= x"000000000000E000";
--                        for i in 13 to 15 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000010000" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"000000000001C000";
--                        for i in 14 to 16 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000010001" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000000038000";
--                        for i in 15 to 17 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000010010" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000000070000";
--                        for i in 16 to 18 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000010011" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"00000000000E0000";
--                        for i in 17 to 19 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000010100" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"00000000001C0000";
--                        for i in 18 to 20 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000010101" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000000380000";
--                        for i in 19 to 21 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000010110" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000000700000";
--                        for i in 20 to 22 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000010111" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000000E00000";
--                        for i in 21 to 23 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000011000" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000001C00000";
--                        for i in 22 to 24 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000011001" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000003800000";
--                        for i in 23 to 25 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000011010" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000007000000";
--                        for i in 24 to 26 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000011011" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"000000000E000000";
--                        for i in 25 to 27 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000011100" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"000000001C000000";
--                        for i in 26 to 28 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000011101" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000038000000";
--                        for i in 27 to 29 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000011110" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000070000000";
--                        for i in 28 to 30 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000011111" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"00000000E0000000";
--                        for i in 29 to 31 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000100000" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"00000001C0000000";
--                        for i in 30 to 32 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000100001" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000380000000";
--                        for i in 31 to 33 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000100010" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000700000000";
--                        for i in 32 to 34 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000100011" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000E00000000";
--                        for i in 33 to 35 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000100100" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000001C00000000";
--                        for i in 34 to 36 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000100101" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000380000000";
--                        for i in 35 to 37 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000100110" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000007000000000";
--                        for i in 36 to 38 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000100111" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"000000E000000000";
--                        for i in 37 to 39 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000101000" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"000001C000000000";
--                        for i in 38 to 40 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000101001" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000038000000000";
--                        for i in 39 to 41 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000101010" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000070000000000";
--                        for i in 40 to 42 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000101011" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"00000E0000000000";
--                        for i in 41 to 43 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000101100" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"00001C0000000000";
--                        for i in 42 to 44 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000101101" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000380000000000";
--                        for i in 43 to 45 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000101110" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000700000000000";
--                        for i in 44 to 46 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000101111" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000E00000000000";
--                        for i in 45 to 47 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000110000" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0001C00000000000";
--                        for i in 46 to 48 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000110001" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0003800000000000";
--                        for i in 47 to 49 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000110010" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0007000000000000";
--                        for i in 48 to 50 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000110011" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"000E000000000000";
--                        for i in 49 to 51 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000110100" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"001C000000000000";
--                        for i in 50 to 52 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000110101" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0038000000000000";
--                        for i in 51 to 53 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000110110" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0070000000000000";
--                        for i in 52 to 54 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000110111" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"00E0000000000000";
--                        for i in 53 to 55 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000111000" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"01C0000000000000";
--                        for i in 54 to 56 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000111001" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0380000000000000";
--                        for i in 55 to 57 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000111010" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0700000000000000";
--                        for i in 56 to 58 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000111011" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0E00000000000000";
--                        for i in 57 to 59 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000111100" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"1C00000000000000";
--                        for i in 58 to 60 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000111101" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"3800000000000000";
--                        for i in 59 to 61 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000111110" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"7000000000000000";
--                        for i in 60 to 62 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"000111111" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"E000000000000000";
--                        for i in 61 to 63 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"001000000" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"C000000000000000";
--                        for i in 62 to 63 loop
--                            assign(i) <= pixel_right;
--                        end loop;
--                    elsif x_column = b"001000001" then
--                        enable_write_l <= '0';
--                        enable_write_r <= x"8000000000000000";
--                        assign(63) <= pixel_right;
--                    else
--                        enable_write_l <= '0';
--                        enable_write_r <= x"0000000000000000";
--                        for i in 0 to D - 1 loop
--                            assign(i) <= (others => '0');
--                        end loop;
--                end if;
    end process assign_process; 

	
	clk_generator_process : process 
	begin
		clk <= not clk;
		wait for 50 ns;
		
		clk <= not clk;
		wait for 50 ns;
	end process clk_generator_process;
	
	
end arquitectura; 